LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY esteira IS
	PORT(PESO: IN BIT;
			BALANCA: IN BIT;
		SERVO_POSITION: OUT BIT_VECTOR (1 DOWNTO 0);--PINO DA POSICAO DO SERVO É : A13 B13
		ESTERIA_ACTIVE:OUT BIT);--PINO ATIVAR ESTEIRA É :A14

end esteira;


ARCHITECTURE esteira_arq OF esteira IS

BEGIN
		PROCESS (PESO,BALANCA)
			BEGIN
				IF BALANCA='1' THEN
					ESTERIA_ACTIVE<='0';
					IF PESO='0' THEN
						SERVO_POSITION<="10";
					ELSIF PESO='1' THEN
						SERVO_POSITION<="01";
					END IF;
				ELSIF BALANCA='0' THEN
					ESTERIA_ACTIVE<='1';
				END IF;
			END PROCESS;
		--SERVO_POSITION<= "10" WHEN PESO='1' ELSE
		--					  "01" WHEN PESO='0';
		--ESTERIA_ACTIVE<= '1' WHEN BALANCA='0' ELSE
			--					'0' WHEN BALANCA='1';
END esteira_arq;
							  